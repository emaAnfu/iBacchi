CIRCUIT C:\Users\aless\Desktop\CarryInverterV2\CarryInverterV2.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* Generators for phi and notCarry
Vin IN 0 PULSE(0 1.2 125p 10p 10p 250p 500p)
*
* MOS devices
MN1 OUT IN 0 0 N1  W= 0.6U L= 0.12U
MP1 OUT IN 1 1 P1  W= 1.8U L= 0.12U
*
*
* Output capacitance
Cadd OUT 0 100fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=1 VTO=0.40 UO=600.000 TOX= 2.0E-9
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=1 VTO=-0.45 UO=200.000 TOX= 2.0E-9
*
* Transient analysis
*
.TEMP 27.0
.tran 0 0.65n 0 1p
.PROBE
.END
