* D:\INGEGNERIA\Microelectronics\iBacchi\Microelectronics Mod. B - Valle\nMOSCaratt\nMosCaratt.sch

* Schematics Version 9.1 - Web Update 1
* Fri Jul 07 09:56:25 2017



** Analysis setup **
.DC LIN V_Vgs 0 3.3 0.01 
.OP 
.LIB "D:\INGEGNERIA\Microelectronics\VALLE\nMOSCaratt\nMosCaratt.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"
.lib "C:\Program Files\OrCAD_Demo\Capture\Library\Pspice\uwind.lib"

.INC "nMosCaratt.net"
.INC "nMosCaratt.als"


.probe


.END
