* D:\INGEGNERIA\Microelectronics\iBacchi\Microelectronics Mod. B - Valle\nMOSCaratt\nMosR0.sch

* Schematics Version 9.1 - Web Update 1
* Fri Jul 07 14:41:11 2017



** Analysis setup **
.DC LIN V_Vds 0 3.3 0.01 
.OP 
.LIB "D:\INGEGNERIA\Microelectronics\VALLE\nMOSCaratt\nMosCaratt.lib"
.LIB "D:\INGEGNERIA\Microelectronics\iBacchi\Microelectronics Mod. B - Valle\nMOSCaratt\nMosCaratt.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"
.lib "C:\Program Files\OrCAD_Demo\Capture\Library\Pspice\uwind.lib"

.INC "nMosR0.net"
.INC "nMosR0.als"


.probe


.END
