* D:\INGEGNERIA\Microelectronics\VALLE\nMOSCaratt\nMosCaratt.sch

* Schematics Version 9.1 - Web Update 1
* Thu Jul 06 11:18:06 2017



** Analysis setup **
.DC LIN V_Vds 0 3.3 0.01 
.OP 
.LIB "D:\INGEGNERIA\Microelectronics\VALLE\nMOSCaratt\nMosCaratt.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"
.lib "C:\Program Files\OrCAD_Demo\Capture\Library\Pspice\uwind.lib"

.INC "nMosCaratt.net"
.INC "nMosCaratt.als"


.probe


.END
